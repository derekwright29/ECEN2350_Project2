module stateMachine();
endmodule
