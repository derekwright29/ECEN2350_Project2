module BCD(count, display);
	input [9:0] count;
	output reg [20:0] display;
	
	
	endmodule